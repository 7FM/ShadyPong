`ifndef CONFIG_SV
`define CONFIG_SV

//`define VGA_640_350_70_Hz
//`define VGA_640_350_85_Hz
//`define VGA_640_400_70_Hz
//`define VGA_640_400_85_Hz
//`define VGA_640_480_60_Hz
//`define VGA_640_480_73_Hz
`define VGA_640_480_75_Hz
//`define VGA_640_480_85_Hz
//`define VGA_640_480_100_Hz
//`define VGA_720_400_85_Hz
//`define VGA_768_576_60_Hz
//`define VGA_768_576_72_Hz
//`define VGA_768_576_75_Hz
//`define VGA_800_600_56_Hz
//`define VGA_800_600_60_Hz
//`define VGA_1024_768_43_Hz_INTERLACED

`endif
